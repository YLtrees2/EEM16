// Code your design here
`include "dassign1.v"