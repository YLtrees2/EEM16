// Code your testbench here
// or browse Examples
`include "dassign1.tb.v"